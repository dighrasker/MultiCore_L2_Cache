module MSHR #() (



);





endmodule